# pat .... like STL file format, user can define the virtual transaction model to replay the bus transaction function
