// define your assertions here ....

