

module dut_dummy( input clock, input reset);

endmodule
