// record TRX to database
